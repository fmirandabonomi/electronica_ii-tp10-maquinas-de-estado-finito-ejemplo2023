library IEEE;
use IEEE.std_logic_1164.all;

entity receptor_ir_tb is
    -- Vacío
end receptor_ir_tb;

architecture tb of receptor_ir_tb is
    -- Declaraciones
begin
    -- Implementación
end architecture;